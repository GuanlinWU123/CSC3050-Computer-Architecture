`timescale 1ns/1ps
`define assert(signal, value) \
        if (signal !== value) begin \
            $display("ASSERTION FAILED in %m: signal != value"); \
            $finish; \
        end

module alu_test;

reg[31:0] instruction, reg_A, reg_B;
wire[31:0] result;
wire[2:0] flags;
alu testalu(instruction, reg_A, reg_B, result, flags);

initial
    begin
    $display("result: ");
    $monitor("%b : %b", testalu.result, testalu.flags);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0000; //add
    reg_A<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
    reg_B<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b1000_0000_0000_0000_0000_0000_0000_0010);
    #10 `assert(testalu.flags, 3'b001);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0001; //addu
    reg_A<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    reg_B<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b1000_0000_0000_0000_0000_0000_0000_0000);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0010; //sub
    reg_A<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    reg_B<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    #10 `assert(testalu.result, 32'b1111_1111_1111_1111_1111_1111_1111_1110);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0011; //subu
    reg_A<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    reg_B<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    #10 `assert(testalu.result, 32'b0111_1111_1111_1111_1111_1111_1111_1110);   

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0100; //and
    reg_A<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    reg_B<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 `assert(testalu.result, 32'b0100_0000_0100_0000_0100_0000_0100_0000);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0111; //nor
    reg_A<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    reg_B<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 `assert(testalu.result, 32'b0010_0010_0010_0010_0010_0010_0010_0010);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0101; //or
    reg_A<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    reg_B<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 `assert(testalu.result, 32'b1101_1101_1101_1101_1101_1101_1101_1101);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_0110; //xor
    reg_A<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    reg_B<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 `assert(testalu.result, 32'b1001_1101_1001_1101_1001_1101_1001_1101);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_1010; //slt
    reg_A<=32'b1000_0000_0000_0000_0000_0000_0000_0011;
    reg_B<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b0000_0000_0000_0000_0000_0000_0000_0001);
    #10 `assert(testalu.flags, 3'b010);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0010_1011; //sltu
    reg_A<=32'b1000_0000_0000_0000_0000_0000_0000_0011;
    reg_B<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 0);
    #10 `assert(testalu.flags, 3'b0);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_1000_0000; //sll
    reg_A<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    reg_B<=32'b1100_0000_0000_0000_0000_0000_0000_0011;
    #10 `assert(testalu.result, 32'b0000_0000_0000_0000_0000_0000_0000_1100);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_1000_0100; //sllv
    reg_A<=32'b0000_0000_0000_0000_0000_0000_0000_1000;
    reg_B<=32'b1100_0000_0000_0000_0000_0000_0000_0011;
    #10 `assert(testalu.result, 32'b00000000000000000000001100000000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_1000_0010; //srl
    reg_A<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    reg_B<=32'b1100_0000_0000_0000_0000_0000_0000_0011;
    #10 `assert(testalu.result, 32'b001100_0000_0000_0000_0000_0000_0000_00);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_1000_0110; //srlv
    reg_A<=32'b0000_0000_0000_0000_0000_0000_0000_1000;
    reg_B<=32'b1100_0000_0000_0000_0000_0000_0000_0011;
    #10 `assert(testalu.result, 32'b0000_0000_1100_0000_0000_0000_0000_0000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0100_0000_0011; //sra
    reg_A<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    reg_B<=32'b1100_0000_0000_0000_0000_0000_0000_0011;
    #10 `assert(testalu.result, 32'b1111_1111_1111_1111_1100_0000_0000_0000);

    #10 instruction<=32'b0000_0000_0000_0001_0000_0000_0000_0111; //srav
    reg_A<=32'b0100_0000_0000_0000_0000_0000_0000_1000;
    reg_B<=32'b0100_0000_0000_0000_0000_0000_0000_0011;
    #10 `assert(testalu.result, 32'b0);

    #10 instruction<=32'b0010_0000_0000_0001_0000_0000_0000_0001; //addi
    reg_A<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    reg_B<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 `assert(testalu.result, 32'b0000_0000_0000_0000_0000_0000_0000_0000);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0010_0100_0000_0001_0000_0000_0000_0001; //addiu
    reg_A<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    reg_B<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 `assert(testalu.result, 32'b0);
    #10 `assert(testalu.flags, 3'b0);

    #10 instruction<=32'b0001_0000_0000_0001_0000_0000_0000_0001; //beq
    reg_A<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    reg_B<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b0000_0000_0000_0000_0000_0000_0000_0000);
    #10 `assert(testalu.flags, 3'b100);

    #10 instruction<=32'b0001_0100_0000_0001_0000_0000_0000_0001; //bne
    reg_A<=32'b1011_1111_1111_1111_1111_1111_1111_1111;
    reg_B<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b1100_0000_0000_0000_0000_0000_0000_0000);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b1000_1100_0000_0001_0000_0000_0000_0001; //lw
    reg_A<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    reg_B<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b1101_1101_1101_1101_1101_1101_1101_1110);
    #10 `assert(testalu.flags, 3'b000);

    #10 instruction<=32'b0010_1000_0000_0001_0000_0000_0000_0010; //slti
    reg_A<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    reg_B<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b0000_0000_0000_0000_0000_0000_0000_0001);
    #10 `assert(testalu.flags, 3'b010);

    #10 instruction<=32'b0010_1100_0000_0001_1000_0000_0000_0001; //sltiu
    reg_A<=32'b0000_0000_0000_0000_1100_0000_0000_0000;
    reg_B<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
    #10 `assert(testalu.result, 32'b0);
    #10 `assert(testalu.flags, 3'b0);

    #10 $finish;
    end
endmodule